module MUX2X1(a0,a1,s,y);
    input a0,a1,s;
    output y;
    not n1(s_n,s);
    and and1(and_1,s_n,a0);
    and and2(and_2,s,a1);
    or or1(y,and_1,and_2);
endmodule
module DEC5T32E(i,en,y);
    input [4:0] i;
    input en;
    output [31:0]y;
    wire in[4:0];
    not(in[0],i[0]);
    not(in[1],i[1]);
    not(in[2],i[2]);
    not(in[3],i[3]);
    not(in[4],i[4]);
    and a0 (y[0],in[0],in[1],in[2],in[3],in[4],en);
    and a1 (y[1],i[0],in[1],in[2],in[3],in[4],en);
    and a2 (y[2],in[0],i[1],in[2],in[3],in[4],en);
    and a3 (y[3],i[0],i[1],in[2],in[3],in[4],en);
    and a4 (y[4],in[0],in[1],i[2],in[3],in[4],en);
    and a5 (y[5],i[0],in[1],i[2],in[3],in[4],en);
    and a6 (y[6],in[0],i[1],i[2],in[3],in[4],en);
    and a7 (y[7],i[0],i[1],i[2],in[3],in[4],en);
    and a8 (y[8],in[0],in[1],in[2],i[3],in[4],en);
    and a9 (y[9],i[0],in[1],in[2],i[3],in[4],en);
    and a10 (y[10],in[0],i[1],in[2],i[3],in[4],en);
    and a11 (y[11],i[0],i[1],in[2],i[3],in[4],en);
    and a12 (y[12],in[0],in[1],i[2],i[3],in[4],en);
    and a13 (y[13],i[0],in[1],i[2],i[3],in[4],en);
    and a14 (y[14],in[0],i[1],i[2],i[3],in[4],en);
    and a15 (y[15],i[0],i[1],i[2],i[3],in[4],en);
    and a16 (y[16],in[0],in[1],in[2],in[3],i[4],en);
    and a17 (y[17],i[0],in[1],in[2],in[3],i[4],en);
    and a18 (y[18],in[0],i[1],in[2],in[3],i[4],en);
    and a19 (y[19],i[0],i[1],in[2],in[3],i[4],en);
    and a20 (y[20],in[0],in[1],i[2],in[3],i[4],en);
    and a21 (y[21],i[0],in[1],i[2],in[3],i[4],en);
    and a22 (y[22],in[0],i[1],i[2],in[3],i[4],en);
    and a23 (y[23],i[0],i[1],i[2],in[3],i[4],en);
    and a24 (y[24],in[0],in[1],in[2],i[3],i[4],en);
    and a25 (y[25],i[0],in[1],in[2],i[3],i[4],en);
    and a26 (y[26],in[0],i[1],in[2],i[3],i[4],en);
    and a27 (y[27],i[0],i[1],in[2],i[3],i[4],en);
    and a28 (y[28],in[0],in[1],i[2],i[3],i[4],en);
    and a29 (y[29],i[0],in[1],i[2],i[3],i[4],en);
    and a30 (y[30],in[0],i[1],i[2],i[3],i[4],en);
    and a31 (y[31],i[0],i[1],i[2],i[3],i[4],en);
endmodule

module MUX32X1(s,en,a31,a30,a29,a28,a27,a26,a25,a24,a23,a22,a21,a20,a19,a18,a17,a16,a15,a14,a13,a12,a11,a10,a9,a8,a7,a6,a5,a4,a3,a2,a1,a0,y);
    input [31:0]s;
    input en;
    input a31,a30,a29,a28,a27,a26,a25,a24,a23,a22,a21,a20,a19,a18,a17,a16,a15,a14,a13,a12,a11,a10,a9,a8,a7,a6,a5,a4,a3,a2,a1,a0;
    output y;
    and and31 (d31,a31,s[31],en);
    and and30 (d30,a30,s[30],en);
    and and29 (d29,a29,s[29],en);
    and and28 (d28,a28,s[28],en);
    and and27 (d27,a27,s[27],en);
    and and26 (d26,a26,s[26],en);
    and and25 (d25,a25,s[25],en);
    and and24 (d24,a24,s[24],en);
    and and23 (d23,a23,s[23],en);
    and and22 (d22,a22,s[22],en);
    and and21 (d21,a21,s[21],en);
    and and20 (d20,a20,s[20],en);
    and and19 (d19,a19,s[19],en);
    and and18 (d18,a18,s[18],en);
    and and17 (d17,a17,s[17],en);
    and and16 (d16,a16,s[16],en);
    and and15 (d15,a15,s[15],en);
    and and14 (d14,a14,s[14],en);
    and and13 (d13,a13,s[13],en);
    and and12 (d12,a12,s[12],en);
    and and11 (d11,a11,s[11],en);
    and and10 (d10,a10,s[10],en);
    and and9 (d9,a9,s[9],en);
    and and8 (d8,a8,s[8],en);
    and and7 (d7,a7,s[7],en);
    and and6 (d6,a6,s[6],en);
    and and5 (d5,a5,s[5],en);
    and and4 (d4,a4,s[4],en);
    and and3 (d3,a3,s[3],en);
    and and2 (d2,a2,s[2],en);
    and and1 (d1,a1,s[1],en);
    and and0 (d0,a0,s[0],en);
    or (y,d0,d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31);
endmodule 

module MUX32X32(a0,a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15,a16,a17,a18,a19,a20,a21,a22,a23,a24,a25,a26,a27,a28,a29,a30,a31,s,y);
    input [31:0]a0,a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15,a16,a17,a18,a19,a20,a21,a22,a23,a24,a25,a26,a27,a28,a29,a30,a31;
    input [4:0]s;
    output [31:0]y;
    wire [31:0] sw;
    DEC5T32E s1(s,1,sw);
    MUX32X1 m0(a0[0]);
endmodule

module D_Latch(D,En,Q,Qn);
    input D,En;
    output Q,Qn;
    wire Sn,Rn,Dn;
    not i0(Dn,D);
    nand i1(Sn,D,En);
    nand i2(Rn,En,Dn);
    nand i3(Q,Sn,Qn);
    nand i4(Qn,Q,Rn);
endmodule

module D_FF(D,Clk,Q,Qn);
    input D,Clk;
    output Q,Qn;
    wire Clkn,Q0,Qn0;
    not i0(Clkn,Clk);
    D_Latch d0(D,Clkn,Q0,Qn0);
    D_Latch d1(Q0,Clk,Q,Qn);
endmodule

module D_FFEC(D,Clk,En,Clrn,Q,Qn);
    input D,Clk,En,Clrn;
    output Q,Qn;
    wire Y0,Y_C;
    MUX2X1 m0(Q,D,En,Y0);
    and i0(Y_C,Y0,Clrn);//and or nand?
    D_FF d0(Y_C,Clk,Q,Qn);
endmodule

module D_FFEC32(D,Clk,En,Clrn,Q,Qn);
    input [31:0] D;
    input Clk,En,Clrn;
    output [31:0] Q,Qn;
    D_FFEC d0 (D[0],Clk,En,Clrn,Q[0],Qn);
    D_FFEC d1 (D[1],Clk,En,Clrn,Q[1],Qn);
    D_FFEC d2 (D[2],Clk,En,Clrn,Q[2],Qn);
    D_FFEC d3 (D[3],Clk,En,Clrn,Q[3],Qn);
    D_FFEC d4 (D[4],Clk,En,Clrn,Q[4],Qn);
    D_FFEC d5 (D[5],Clk,En,Clrn,Q[5],Qn);
    D_FFEC d6 (D[6],Clk,En,Clrn,Q[6],Qn);
    D_FFEC d7 (D[7],Clk,En,Clrn,Q[7],Qn);
    D_FFEC d8 (D[8],Clk,En,Clrn,Q[8],Qn);
    D_FFEC d9 (D[9],Clk,En,Clrn,Q[9],Qn);
    D_FFEC d10 (D[10],Clk,En,Clrn,Q[10],Qn);
    D_FFEC d11 (D[11],Clk,En,Clrn,Q[11],Qn);
    D_FFEC d12 (D[12],Clk,En,Clrn,Q[12],Qn);
    D_FFEC d13 (D[13],Clk,En,Clrn,Q[13],Qn);
    D_FFEC d14 (D[14],Clk,En,Clrn,Q[14],Qn);
    D_FFEC d15 (D[15],Clk,En,Clrn,Q[15],Qn);
    D_FFEC d16 (D[16],Clk,En,Clrn,Q[16],Qn);
    D_FFEC d17 (D[17],Clk,En,Clrn,Q[17],Qn);
    D_FFEC d18 (D[18],Clk,En,Clrn,Q[18],Qn);
    D_FFEC d19 (D[19],Clk,En,Clrn,Q[19],Qn);
    D_FFEC d20 (D[20],Clk,En,Clrn,Q[20],Qn);
    D_FFEC d21 (D[21],Clk,En,Clrn,Q[21],Qn);
    D_FFEC d22 (D[22],Clk,En,Clrn,Q[22],Qn);
    D_FFEC d23 (D[23],Clk,En,Clrn,Q[23],Qn);
    D_FFEC d24 (D[24],Clk,En,Clrn,Q[24],Qn);
    D_FFEC d25 (D[25],Clk,En,Clrn,Q[25],Qn);
    D_FFEC d26 (D[26],Clk,En,Clrn,Q[26],Qn);
    D_FFEC d27 (D[27],Clk,En,Clrn,Q[27],Qn);
    D_FFEC d28 (D[28],Clk,En,Clrn,Q[28],Qn);
    D_FFEC d29 (D[29],Clk,En,Clrn,Q[29],Qn);
    D_FFEC d30 (D[30],Clk,En,Clrn,Q[30],Qn);
    D_FFEC d31 (D[31],Clk,En,Clrn,Q[31],Qn);
endmodule

module REG32(D,En,Clk,Clrn,Q31,Q30,Q29,Q28,Q27,Q26,Q25,Q24,Q23,Q22,Q21,Q20,Q19,Q18,Q17,Q16,Q15,Q14,Q13,Q12,Q11,Q10,Q9,Q8,Q7,Q6,Q5,Q4,Q3,Q2,Q1,Q0);
    input [31:0]D,En;
    input Clk,Clrn;
    output [31:0] Q31,Q30,Q29,Q28,Q27,Q26,Q25,Q24,Q23,Q22,Q21,Q20,Q19,Q18,Q17,Q16,Q15,Q14,Q13,Q12,Q11,Q10,Q9,Q8,Q7,Q6,Q5,Q4,Q3,Q2,Q1,Q0;
    D_FFEC32 q31 (D,Clk,En[31],Clrn,Q31);
    D_FFEC32 q30 (D,Clk,En[30],Clrn,Q30);
    D_FFEC32 q29 (D,Clk,En[29],Clrn,Q29);
    D_FFEC32 q28 (D,Clk,En[28],Clrn,Q28);
    D_FFEC32 q27 (D,Clk,En[27],Clrn,Q27);
    D_FFEC32 q26 (D,Clk,En[26],Clrn,Q26);
    D_FFEC32 q25 (D,Clk,En[25],Clrn,Q25);
    D_FFEC32 q24 (D,Clk,En[24],Clrn,Q24);
    D_FFEC32 q23 (D,Clk,En[23],Clrn,Q23);
    D_FFEC32 q22 (D,Clk,En[22],Clrn,Q22);
    D_FFEC32 q21 (D,Clk,En[21],Clrn,Q21);
    D_FFEC32 q20 (D,Clk,En[20],Clrn,Q20);
    D_FFEC32 q19 (D,Clk,En[19],Clrn,Q19);
    D_FFEC32 q18 (D,Clk,En[18],Clrn,Q18);
    D_FFEC32 q17 (D,Clk,En[17],Clrn,Q17);
    D_FFEC32 q16 (D,Clk,En[16],Clrn,Q16);
    D_FFEC32 q15 (D,Clk,En[15],Clrn,Q15);
    D_FFEC32 q14 (D,Clk,En[14],Clrn,Q14);
    D_FFEC32 q13 (D,Clk,En[13],Clrn,Q13);
    D_FFEC32 q12 (D,Clk,En[12],Clrn,Q12);
    D_FFEC32 q11 (D,Clk,En[11],Clrn,Q11);
    D_FFEC32 q10 (D,Clk,En[10],Clrn,Q10);
    D_FFEC32 q9 (D,Clk,En[9],Clrn,Q9);
    D_FFEC32 q8 (D,Clk,En[8],Clrn,Q8);
    D_FFEC32 q7 (D,Clk,En[7],Clrn,Q7);
    D_FFEC32 q6 (D,Clk,En[6],Clrn,Q6);
    D_FFEC32 q5 (D,Clk,En[5],Clrn,Q5);
    D_FFEC32 q4 (D,Clk,En[4],Clrn,Q4);
    D_FFEC32 q3 (D,Clk,En[3],Clrn,Q3);
    D_FFEC32 q2 (D,Clk,En[2],Clrn,Q2);
    D_FFEC32 q1 (D,Clk,En[1],Clrn,Q1);
    D_FFEC32 q0 (D,Clk,En[0],Clrn,Q0);
    assign Q0 = 0;
endmodule

module REGFILE(Ra,Rb,D,Wr,We,Clk,Clrn,Qa,Qb);
    input [4:0] Ra,Rb,Wr;
    input [31:0] D;
    input We,Clk,Clrn;
    output [31:0]Qa,Qb;
    wire [31:0] Y_mux,Q31_reg32,Q30_reg32,Q29_reg32,Q28_reg32,Q27_reg32,Q26_reg32,Q25_reg32,Q24_reg32,Q23_reg32,Q22_reg32,Q21_reg32,Q20_reg32,Q19_reg32,Q18_reg32,Q17_reg32,Q16_reg32,Q15_reg32,Q14_reg32,Q13_reg32,Q12_reg32,Q11_reg32,Q10_reg32,Q9_reg32,Q8_reg32,Q7_reg32,Q6_reg32,Q5_reg32,Q4_reg32,Q3_reg32,Q2_reg32,Q1_reg32,Q0_reg32;
    DEC5T32E dec(Wr,We,Y_mux);
    REG32 r1 (D,Y_mux,Clk,Clrn,Q31_reg32,Q30_reg32,Q29_reg32,Q28_reg32,Q27_reg32,Q26_reg32,Q25_reg32,Q24_reg32,Q23_reg32,Q22_reg32,Q21_reg32,Q20_reg32,Q19_reg32,Q18_reg32,Q17_reg32,Q16_reg32,Q15_reg32,Q14_reg32,Q13_reg32,Q12_reg32,Q11_reg32,Q10_reg32,Q9_reg32,Q8_reg32,Q7_reg32,Q6_reg32,Q5_reg32,Q4_reg32,Q3_reg32,Q2_reg32,Q1_reg32,Q0_reg32);
    MUX32X32 select1();
    MUX32X32 select2();
endmodule