module DEC2T4E(i0,i1,en,y0,y1,y2,y3);
    input i0,i1,en;
    output y0,y1,y2,y3;
    assign y0 = (~i0)&(~i1)&en;
    assign y1 = (~i0)&i1&en;
    assign y2 = i0&(~i1)&en;
    assign y3 = i0&i1&en;
endmodule

module DEC5T32E(i,en,y);
    input [4:0]i;
    input en;
    output [31:0]y;
    function [31:0]dec;
        input [31:0]i;
        output [31:0]y;
        case (i)
            2'b00000:dec = 00000000000000000000000000000001;
            2'b00001:dec = 00000000000000000000000000000010;
            2'b00010:dec = 00000000000000000000000000000100;
            2'b00011:dec = 00000000000000000000000000001000;
            2'b00100:dec = 00000000000000000000000000010000;
            2'b00101:dec = 00000000000000000000000000100000;
            2'b00110:dec = 00000000000000000000000001000000;
            2'b00111:dec = 00000000000000000000000010000000;
            2'b01000:dec = 00000000000000000000000100000000;
            2'b01001:dec = 00000000000000000000001000000000;
            2'b01010:dec = 00000000000000000000010000000000;
            2'b01011:dec = 00000000000000000000100000000000;
            2'b01100:dec = 00000000000000000001000000000000;
            2'b01101:dec = 00000000000000000010000000000000;
            2'b01110:dec = 00000000000000000100000000000000;
            2'b01111:dec = 00000000000000001000000000000000;
            2'b10000:dec = 00000000000000010000000000000000;
            2'b10001:dec = 00000000000000100000000000000000;
            2'b10010:dec = 00000000000001000000000000000000;
            2'b10011:dec = 00000000000010000000000000000000;
            2'b10100:dec = 00000000000100000000000000000000;
            2'b10101:dec = 00000000001000000000000000000000;
            2'b10110:dec = 00000000010000000000000000000000;
            2'b10111:dec = 00000000100000000000000000000000;
            2'b11000:dec = 00000001000000000000000000000000;
            2'b11001:dec = 00000010000000000000000000000000;
            2'b11010:dec = 00000100000000000000000000000000;
            2'b11011:dec = 00001000000000000000000000000000;
            2'b11100:dec = 00010000000000000000000000000000;
            2'b11101:dec = 00100000000000000000000000000000;
            2'b11110:dec = 01000000000000000000000000000000;
            2'b11111:dec = 10000000000000000000000000000000;
        endcase
    assign y = dec(i);
    if (en==2'b0)) begin
        assign y = 2'b00000000000000000000000000000000;  
    end
endmodule